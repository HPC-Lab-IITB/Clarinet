// Copyright (c) 2016-2020 Bluespec, Inc. All Rights Reserved

package CPU_Stage2;

// ================================================================
// This is Stage 2 of the CPU.
// It is the "DM" stage ("Data Memory"), which is the main function.

// However, this stage also contains all other (potentially) long-latency
// operations:
//    MBox ("M" extension ops, integer multiply/divide)
//    FDBox ("FD" extension ops, single and double precision floating point)

// This stage sends out Tandem Verifier information for pipelined instructions

// Note: $displays are indented by (stage num x 4) spaces.
// for traditional pipeline display
//     IF
//         DM
//             WB
// i.e., 8 spaces for this stage.

// ================================================================
// Exports

export
CPU_Stage2_IFC (..),
mkCPU_Stage2;

// ================================================================
// BSV library imports

import FIFOF        :: *;
import GetPut       :: *;
import ClientServer :: *;
import ConfigReg    :: *;

// ----------------
// BSV additional libs

import Cur_Cycle  :: *;

// ================================================================
// Project imports

import ISA_Decls     :: *;

import TV_Info       :: *;

import CPU_Globals   :: *;
import Near_Mem_IFC  :: *;
import CSR_RegFile   :: *;    // For SATP, SSTATUS, MSTATUS

`ifdef SHIFT_SERIAL
import Shifter_Box  :: *;
`endif

`ifdef ISA_M
import RISCV_MBox  :: *;
`endif

`ifdef ISA_F
import FBox_Top    :: *;
import FBox_Core   :: *;   // For fv_nanbox function
`endif

`ifdef ROCC               //Stage 2 dispatches to PositAccel
import PositAccel      :: *;
`endif

`ifdef ACCEL               //Stage 2 dispatches to PositAccel
import PositAccel      :: *;
`endif
// ================================================================
// Interface

interface CPU_Stage2_IFC;
   // ---- Reset
   interface Server #(Token, Token) server_reset;

   // ---- Output
   (* always_ready *)
   method Output_Stage2  out;

   (* always_ready *)
   method Action deq;

   // ---- Input
   (* always_ready *)
   method Action enq (Data_Stage1_to_Stage2 x);

   (* always_ready *)
   method Action set_full (Bool full);
endinterface

// ================================================================
// Implementation module

module mkCPU_Stage2 #(Bit #(4)         verbosity,
		      CSR_RegFile_IFC  csr_regfile,    // for SATP and SSTATUS: TODO carry in Data_Stage1_to_Stage2
		      DMem_IFC         dcache)
                    (CPU_Stage2_IFC);

   FIFOF #(Token) f_reset_reqs <- mkFIFOF;
   FIFOF #(Token) f_reset_rsps <- mkFIFOF;

   Reg #(Bool)                  rg_resetting  <- mkReg (False);
   Reg #(Bool)                  rg_full       <- mkReg (False);
   Reg #(Data_Stage1_to_Stage2) rg_stage2     <- mkRegU;    // From Stage 1

   // ----------------
   // Serial shifter box

`ifdef SHIFT_SERIAL
   Shifter_Box_IFC shifter_box <- mkShifter_Box;
`endif

   // ----------------
   // Integer multiply/divide box

`ifdef ISA_M
   RISCV_MBox_IFC mbox <- mkRISCV_MBox;
`endif

   // ----------------
   // Floating point box

`ifdef ISA_F
   FBox_Top_IFC fbox <- mkFBox_Top (0);
`endif
  // ----------------
   // PositAccel Wrapper

`ifdef ROCC//instantiate the wrapper PositAccel
   Wrapper_IFC wrap <- mkPositAccel ; 
`endif

`ifdef ACCEL//instantiate the wrapper PositAccel
   Wrapper_IFC wrap <- mkPositAccel ; 
`endif
   // ----------------

   let bypass_base = Bypass {bypass_state: BYPASS_RD_NONE,
			     rd:           rg_stage2.rd,
			     rd_val:       rg_stage2.val1
			     };

`ifdef ISA_F
   let fbypass_base = FBypass {bypass_state: BYPASS_RD_NONE,
			       rd:           rg_stage2.rd,
			       rd_val:       rg_stage2.fval1
			       };

// Bypass logic for the posit RF
`ifdef POSIT
   let pbypass_base = PBypass {bypass_state: BYPASS_RD_NONE,
			       rd:           rg_stage2.rd,
			       rd_val:       rg_stage2.pval1
			       };

`endif
`endif

`ifdef ROCC               //Bypass Logic for ACCEL i.e PositAccel
   let roccbypass_base = roccBypass {bypass_state: BYPASS_RD_NONE,
			       rd:           rg_stage2.rd,
			       rd_val:       rg_stage2.roccval1
			       };
`endif


`ifdef ACCEL               //Bypass Logic for ACCEL i.e PositAccel
   let accelbypass_base = AccelBypass {bypass_state: BYPASS_RD_NONE,
			       rd:           rg_stage2.rd,
			       rd_val:       rg_stage2.accelval1
			       };
`endif

   let data_to_stage3_base = Data_Stage2_to_Stage3 {
        priv:      rg_stage2.priv
      , pc:        rg_stage2.pc
      , instr:     rg_stage2.instr
`ifdef ISA_F
      , rd_in_fpr: False
      , upd_flags: False
      , fpr_flags: 0
      , frd_val  : rg_stage2.fval1
`ifdef POSIT
      , no_rd_upd: False
      , rd_in_ppr: False
      , prd_val  : rg_stage2.pval1
`endif
`endif
      ,	rd_valid:  False
      , rd:        rg_stage2.rd
      , rd_val:    rg_stage2.val1

`ifdef ROCC               //changes maybe required 
      , no_rd_upd: False
      , rd_in_ppr: False
      , prd_val  : rg_stage2.roccval1

`endif

`ifdef ACCEL               //changes maybe required 
      , no_rd_upd: False
      , rd_in_ppr: False
      , prd_val  : rg_stage2.accelval1

`endif
`ifdef INCLUDE_TANDEM_VERIF
      , trace_data: rg_stage2.trace_data
`endif
   };

   let  trap_info_dmem = Trap_Info {epc:      rg_stage2.pc,
				    exc_code: dcache.exc_code,
				    tval:     rg_stage2.addr };

`ifdef ISA_F
   // The FBox can only generate ILLEGAL Instruction exceptions
   let  trap_info_fbox = Trap_Info {epc:      rg_stage2.pc,
				    exc_code: exc_code_ILLEGAL_INSTRUCTION,
				    tval:     0 };
`endif

   // ----------------------------------------------------------------
   // BEHAVIOR

   rule rl_reset_begin;
      f_reset_reqs.deq;
      rg_full <= False;
      rg_resetting <= True;
`ifdef ISA_F
      fbox.server_reset.request.put (?);
`endif
   endrule

   rule rl_reset_end (rg_resetting);
      rg_resetting <= False;

`ifdef ISA_F
      let res <- fbox.server_reset.response.get;
`endif

`ifdef ROCC
       let rocc_resp <-wrap.server_reset.response.get;    //server response when PositAccel is set
`endif



`ifdef ACCEL
       let accel_resp <-wrap.server_reset.response.get;    //server response when PositAccel is set
`endif

      f_reset_rsps.enq (?);
   endrule


 

   // ----------------
   // Combinational output function

   function Output_Stage2 fv_out;
      Output_Stage2 output_stage2 = ?;

      // This stage is empty
      if (! rg_full) begin
	 output_stage2 = Output_Stage2 {ostatus         : OSTATUS_EMPTY,
					trap_info       : ?,
					data_to_stage3  : ?,
					bypass          : no_bypass
`ifdef ISA_F
                                      , fbypass         : no_fbypass

`ifdef POSIT
                                      , pbypass         : no_pbypass

`endif
`endif


`ifdef ROCC
                                      , roccbypass         : no_roccbypass
`endif

`ifdef ACCEL
                                      , accelbypass         : no_accelbypass
`endif

`ifdef INCLUDE_TANDEM_VERIF
	                              , trace_data      : ?
`endif
				       };
      end

      // This stage is just relaying ALU results from previous stage to next stage
      else if (rg_stage2.op_stage2 == OP_Stage2_ALU) begin
	 let data_to_stage3 = data_to_stage3_base;
	 data_to_stage3.rd_valid = True;

	 let bypass = bypass_base;
	 bypass.bypass_state = BYPASS_RD_RDVAL;

	 output_stage2 = Output_Stage2 {ostatus         : OSTATUS_PIPE,
					trap_info       : ?,
					data_to_stage3  : data_to_stage3,
					bypass          : bypass
`ifdef ISA_F
                                      , fbypass         : no_fbypass

`ifdef POSIT
                                      , pbypass         : no_pbypass
`endif
`endif
`ifdef ROCC
                                      , roccbypass         : no_roccbypass
`endif

					};
      end

      // This stage is doing a LOAD or AMO
      else if (   (rg_stage2.op_stage2 == OP_Stage2_LD)
`ifdef ISA_A
	       || (rg_stage2.op_stage2 == OP_Stage2_AMO)
`endif
	       )
	 begin
	    let ostatus = (  (! dcache.valid)
			   ? OSTATUS_BUSY
			   : (  dcache.exc
			      ? OSTATUS_NONPIPE
			      : OSTATUS_PIPE));

	    WordXL result = truncate (dcache.word64);

            let funct3 = instr_funct3 (rg_stage2.instr);

	    let data_to_stage3 = data_to_stage3_base;
	    data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);

`ifdef ISA_F
            data_to_stage3.rd_in_fpr = rg_stage2.rd_in_fpr;
            // A FPR load
            if (rg_stage2.rd_in_fpr) begin
`ifdef ISA_D
               // Both FLW and FLD are legal instructions
               // A FLW result
               if (funct3 == f3_FLW)
                  // needs nan-boxing when destined for a DP register file
                  data_to_stage3.frd_val = fv_nanbox (dcache.word64);

               // A FLD result
               else
                  data_to_stage3.frd_val = dcache.word64;
`else
               // Only FLW is a legal instruction
               data_to_stage3.frd_val = truncate (dcache.word64);
`endif
            end
`ifdef POSIT
            // A PPR load
            else if (rg_stage2.rd_in_ppr) begin
               // Only PLW is a legal instruction
               data_to_stage3.prd_val = truncate (dcache.word64);
            end
            data_to_stage3.rd_in_ppr = rg_stage2.rd_in_ppr;
`endif
`endif
            // GPR loads
	    data_to_stage3.rd_val   = result;


`ifdef ROCC       //need to change
            // A PPR load
             if (rg_stage2.rd_in_ppr) begin
               // Only PLW is a legal instruction
               //It needs to be checked
               data_to_stage3.prd_val = truncate (dcache.word64);
            end
            data_to_stage3.rd_in_ppr = rg_stage2.rd_in_ppr;
`endif

`ifdef ACCEL       //need to change
            // A PPR load
             if (rg_stage2.rd_in_ppr) begin
               // Only PLW is a legal instruction
               //It needs to be checked
               data_to_stage3.prd_val = truncate (dcache.word64);
            end
            data_to_stage3.rd_in_ppr = rg_stage2.rd_in_ppr;
`endif


            // Update the bypass channel, if not trapping (NONPIPE)
	    let bypass = bypass_base;
`ifdef ISA_F
	    let fbypass = fbypass_base;
`ifdef POSIT
	    let pbypass = pbypass_base;
`endif
`endif

`ifdef ROCC
	    let roccbypass = roccbypass_base;
`endif

`ifdef ACCEL
	    let accelbypass = accelbypass_base;
`endif



	    if (ostatus != OSTATUS_NONPIPE) begin
`ifdef ISA_F
               // Bypassing FPR value.
               if (rg_stage2.rd_in_fpr) begin
		  // Choose one of the following two options

		  // Option 1: longer critical path, since the data is bypassed back into previous stage.
		  // We use data_to_stage3.rd_val since nanboxing has been done.
		  // fbypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
		  // fbypass.rd_val       = data_to_stage3.frd_val;

		  // Option 2: shorter critical path, since the data is not bypassed into previous stage,
		  // (the bypassing is effectively delayed until the next stage).
		  fbypass.bypass_state = BYPASS_RD;
               end
`ifdef POSIT
               // Bypassing PPR value.
               else if (rg_stage2.rd_in_ppr) begin
		  // Choose one of the following two options

		  // Option 1: longer critical path, since the data is bypassed back into previous stage.
		  // We use data_to_stage3.rd_val since nanboxing has been done.
		  // pbypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
		  // pbypass.rd_val       = data_to_stage3.prd_val;

		  // Option 2: shorter critical path, since the data is not bypassed into previous stage,
		  // (the bypassing is effectively delayed until the next stage).
		  pbypass.bypass_state = BYPASS_RD;
               end
`endif
`endif


               // Bypassing GPR values
               if (rg_stage2.rd != 0) begin    // TODO: is this test necessary?
		  // Choose one of the following two options

		  // Option 1: longer critical path, since the data is bypassed back into previous stage.
		  // We use data_to_stage3.rd_val since nanboxing has been done.
		  // bypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
		  // bypass.rd_val       = result;

		  // Option 2: shorter critical path, since the data is not bypassed into previous stage,
		  // (the bypassing is effectively delayed until the next stage).
		  bypass.bypass_state = BYPASS_RD;
	       end
	    end


`ifdef ROCC
               // Bypassing PPR value.
               else if (rg_stage2.rd_in_ppr) begin
		  // Choose one of the following two options

		  // Option 1: longer critical path, since the data is bypassed back into previous stage.
		  // We use data_to_stage3.rd_val since nanboxing has been done.
		  // pbypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
		  // pbypass.rd_val       = data_to_stage3.prd_val;

		  // Option 2: shorter critical path, since the data is not bypassed into previous stage,
		  // (the bypassing is effectively delayed until the next stage).
		  roccbypass.bypass_state = BYPASS_RD;
               end
`endif

`ifdef ACCEL
               // Bypassing PPR value.
               else if (rg_stage2.rd_in_ppr) begin
		  // Choose one of the following two options

		  // Option 1: longer critical path, since the data is bypassed back into previous stage.
		  // We use data_to_stage3.rd_val since nanboxing has been done.
		  // pbypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
		  // pbypass.rd_val       = data_to_stage3.prd_val;

		  // Option 2: shorter critical path, since the data is not bypassed into previous stage,
		  // (the bypassing is effectively delayed until the next stage).
		  accelbypass.bypass_state = BYPASS_RD;
               end
`endif


`ifdef INCLUDE_TANDEM_VERIF
	    let trace_data = rg_stage2.trace_data;
`ifdef ISA_F
            if (rg_stage2.rd_in_fpr) begin
               trace_data.word5 = data_to_stage3.frd_val;

               // Update MSTATUS.FS in trace packet
	       let new_mstatus = csr_regfile.mv_update_mstatus_fs (fs_xs_dirty);
               trace_data = fv_trace_update_mstatus_fs (trace_data, new_mstatus);
            end else
`endif
               trace_data.word1 = data_to_stage3.rd_val;

            data_to_stage3.trace_data = trace_data;
`endif

            output_stage2 = Output_Stage2 {ostatus         : ostatus,
					   trap_info       : trap_info_dmem,
					   data_to_stage3  : data_to_stage3,
					   bypass          : bypass
`ifdef ISA_F
                                         , fbypass         : fbypass
`ifdef POSIT
                                         , pbypass         : no_pbypass
`endif
`endif

`ifdef ROCC
                                         , roccbypass         : no_roccbypass
`endif

`ifdef ACCEL
                                         , accelbypass         : no_accelbypass
`endif
`ifdef INCLUDE_TANDEM_VERIF
                                         , trace_data      : trace_data
`endif
					   };
	 end

      // This stage is doing a STORE
      else if (rg_stage2.op_stage2 == OP_Stage2_ST) begin
	 let ostatus = (  (! dcache.valid)
			     ? OSTATUS_BUSY
			     : (  dcache.exc
				? OSTATUS_NONPIPE
				: OSTATUS_PIPE));

	 let data_to_stage3 = data_to_stage3_base;
	 data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);
	 data_to_stage3.rd       = 0;

	 output_stage2 = Output_Stage2 {ostatus         : ostatus,
					trap_info       : trap_info_dmem,
					data_to_stage3  : data_to_stage3,
					bypass          : no_bypass
`ifdef ISA_F
                                      , fbypass         : no_fbypass
`ifdef POSIT
                                      , pbypass         : no_pbypass
`endif
`endif
`ifdef ROCC
                                      , roccbypass         : no_roccbypass
`endif
`ifdef ACCEL
                                      , accelbypass         : no_accelbypass
`endif
`ifdef INCLUDE_TANDEM_VERIF
                                      , trace_data      : trace_data
`endif
					};
      end

`ifdef SHIFT_SERIAL
      // This stage is doing a serial shift
      else if (rg_stage2.op_stage2 == OP_Stage2_SH) begin
	 let ostatus = ((! shifter_box.valid) ? OSTATUS_BUSY : OSTATUS_PIPE);

	 let result = shifter_box.word;

	 let data_to_stage3 = data_to_stage3_base;
	 data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);
	 data_to_stage3.rd_val   = result;

	 let bypass = bypass_base;
	 bypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
	 bypass.rd_val       = result;

`ifdef INCLUDE_TANDEM_VERIF
	 let trace_data            = rg_stage2.trace_data;
	 trace_data.word1          = result;
	 data_to_stage3.trace_data = trace_data;
`endif

	 output_stage2 = Output_Stage2 {ostatus         : ostatus,
					trap_info       : ?,
					data_to_stage3  : data_to_stage3,
					bypass          : bypass
`ifdef ISA_F
                                      , fbypass         : no_fbypass
`ifdef POSIT
                                      , pbypass         : no_pbypass
`endif
`endif
`ifdef ROCC
                                      , roccbypass         : no_roccbypass
`endif

`ifdef INCLUDE_TANDEM_VERIF
                                      , trace_data      : trace_data
`endif
					};
      end
`endif

`ifdef ISA_M
      // This stage is doing an integer multiply/divide
      else if (rg_stage2.op_stage2 == OP_Stage2_M) begin
	 let ostatus = ((! mbox.valid) ? OSTATUS_BUSY : OSTATUS_PIPE);

	 let result = mbox.word;

	 let data_to_stage3 = data_to_stage3_base;
	 data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);
	 data_to_stage3.rd_val   = result;

	 let bypass = bypass_base;
	 bypass.bypass_state = ((ostatus == OSTATUS_PIPE) ? BYPASS_RD_RDVAL : BYPASS_RD);
	 bypass.rd_val       = result;

`ifdef INCLUDE_TANDEM_VERIF
	 let trace_data            = rg_stage2.trace_data;
	 trace_data.word1          = result;
	 data_to_stage3.trace_data = trace_data;
`endif

	 output_stage2 = Output_Stage2 {ostatus         : ostatus,
					trap_info       : ?,
					data_to_stage3  : data_to_stage3,
					bypass          : bypass
`ifdef ISA_F
                                      , fbypass         : no_fbypass
`ifdef POSIT
                                      , pbypass         : no_pbypass
`endif
`endif
`ifdef ROCC
                                      , roccbypass         : no_roccbypass
`endif
`ifdef INCLUDE_TANDEM_VERIF
                                      , trace_data      : trace_data
`endif
					};
      end
`endif

`ifdef ISA_F
      // This stage is doing a floating point op
      else if (rg_stage2.op_stage2 == OP_Stage2_FD) begin
	 let ostatus = ((! fbox.valid) ? OSTATUS_BUSY : OSTATUS_PIPE);

         // Extract fields from FBOX result
	 match {.value, .fflags} = fbox.word;

	 let data_to_stage3      = data_to_stage3_base;
	 data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);
`ifdef ISA_D
	 data_to_stage3.frd_val  = value;
`else
	 data_to_stage3.frd_val  = truncate (value);
`endif
         data_to_stage3.rd_in_fpr= rg_stage2.rd_in_fpr;
         data_to_stage3.upd_flags= True;
         data_to_stage3.fpr_flags= fflags;
`ifdef POSIT
         data_to_stage3.no_rd_upd= rg_stage2.no_rd_upd;
         data_to_stage3.rd_in_prf= rg_stage2.rd_in_prf;
         data_to_stage3.prd_val  = truncate (value);
`endif
`ifdef RV64
         data_to_stage3.rd_val   = value;
`else
         data_to_stage3.rd_val   = truncate (value);
`endif

	 let bypass              = bypass_base;
         let fbypass             = fbypass_base;
`ifdef POSIT
         let pbypass             = pbypass_base;
`endif
         // result is meant for a FPR
         if (rg_stage2.rd_in_fpr) begin
            fbypass.bypass_state    = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
`ifdef ISA_D
            fbypass.rd_val          = value;
`else
            fbypass.rd_val          = truncate (value);
`endif
         end

`ifdef POSIT
         else if ((rg_stage2.rd_in_prf) || (rg_stage2.no_rd_upd)) begin
            if ((rg_stage2.rd_in_prf) && (!rg_stage2.no_rd_upd)) begin
               pbypass.bypass_state = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
               pbypass.rd_val       = truncate (value);
            end
         end
`endif

         // result is meant for a GPR
         else begin
            bypass.bypass_state     = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
`ifdef RV64
            bypass.rd_val           = (value);
`else
            bypass.rd_val           = truncate (value);
`endif
          end

         // -----
`ifdef INCLUDE_TANDEM_VERIF
	 let trace_data = rg_stage2.trace_data;

         if (rg_stage2.rd_in_fpr) begin
            trace_data.word5 = data_to_stage3.frd_val;
         end else begin
            trace_data.word1 = data_to_stage3.rd_val;
         end

	 data_to_stage3.trace_data = trace_data;
 end
`endif

 //--------------------------------------------------------------------
`ifdef ROCC
      // This stage is doing Posit accelerator op
       if (rg_stage2.op_stage2 == OP_Stage2_ROCC) begin  


	     let ostatus = ((! wrap.valid) ? OSTATUS_BUSY : OSTATUS_PIPE); //set status as per posit accel
//instantiation of positaccel has been done using wrap 

    
     // Extract fields from PositAccel result which are necessary to be sent to writeback stage(Stage 3)(clarify this that what all to be sent)

//if xd=0 do not wait for response from wrapper else wait for the response and then proceed

//funct3 in Accelerator is termed as rg_sel-where rg_sel[2] is xd;rg_sel[1] is xs1;rg_sel[0] is xs2.(in terms of RoCC format)
            
          let data_to_stage3  = data_to_stage3_base;
          let  xd  =rg_stage.funct3[2]; //the msb bit of funct3,in RoCC terms its xd
          
	     if((!xd)==0) begin
         Wrapper_in_res rocc_resp=  ff_ROCCRsp.first; //extracting the response from PositAccel in accel_resp
	     data_to_stage3.prd_val  = rocc_resp.result; //accelerator result
         end
         data_to_stage3.no_rd_upd= rg_stage2.no_rd_upd;
	 data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);
         data_to_stage3.rd_in_ppr= rg_stage2.rd_in_ppr;
       
         
	let bypass                = bypass_base;
        let roccbypass           = roccbypass_base;  

         // result is meant for a PPR
         if (rg_stage2.rd_in_ppr) begin
            roccbypass.bypass_state    = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
            roccbypass.rd_val          = value;

         end


         // result is meant for a GPR (while using vector operations)
         else begin
            bypass.bypass_state     = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
`ifdef RV64
            bypass.rd_val           = (value);
`else
            bypass.rd_val           = truncate (value);
`endif
          end
 end
`endif

 // -----------------------------------------------------
//--------------------------------------------------------------------
`ifdef ACCEL
      // This stage is doing Posit accelerator op
       if (rg_stage2.op_stage2 == OP_Stage2_ACCEL) begin  


	     let ostatus = ((! wrap.valid) ? OSTATUS_BUSY : OSTATUS_PIPE); //set status as per posit accel
//instantiation of positaccel has been done using wrap 

    
     // Extract fields from PositAccel result which are necessary to be sent to writeback stage(Stage 3)(clarify this that what all to be sent)

//if xd=0 do not wait for response from wrapper else wait for the response and then proceed

//funct3 in Accelerator is termed as rg_sel-where rg_sel[2] is xd;rg_sel[1] is xs1;rg_sel[0] is xs2.(in terms of RoCC format)
            
          let data_to_stage3  = data_to_stage3_base;
          let  xd  =rg_stage.funct3[2]; //the msb bit of funct3,in RoCC terms its xd
          
	     if((!xd)==0) begin
         Wrapper_in_res accel_resp=  ff_ROCCRsp.first; //extracting the  response from PositAccel in accel_resp
	     data_to_stage3.prd_val  = accel_resp.result; //accelerator result
         end
         data_to_stage3.no_rd_upd= rg_stage2.no_rd_upd;
	 data_to_stage3.rd_valid = (ostatus == OSTATUS_PIPE);
         data_to_stage3.rd_in_ppr= rg_stage2.rd_in_ppr;
       
         
	let bypass                = bypass_base;
        let accelbypass           = accelbypass_base;  

         // result is meant for a PPR
         if (rg_stage2.rd_in_ppr) begin
            accelbypass.bypass_state    = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
            accelbypass.rd_val          = value;

         end


         // result is meant for a GPR (while using vector operations)
         else begin
            bypass.bypass_state     = ((ostatus==OSTATUS_PIPE) ? BYPASS_RD_RDVAL
                                                               : BYPASS_RD);
`ifdef RV64
            bypass.rd_val           = (value);
`else
            bypass.rd_val           = truncate (value);
`endif
          end
 end
`endif

 // -----------------------------------------------------


//stage 2 outputs
	 output_stage2 = Output_Stage2 {ostatus         : ostatus,
					trap_info       : trap_info_fbox,
					data_to_stage3  : data_to_stage3,
					bypass          : bypass
`ifdef ISA_F
                                      , fbypass         : fbypass
`ifdef POSIT
                                      , pbypass         : pbypass
`endif
`endif

`ifdef ROCC
                                      , roccbypass         : roccbypass
`endif

`ifdef ACCEL
                                      , accelbypass         : accelbypass
`endif
`ifdef INCLUDE_TANDEM_VERIF
                                      , trace_data      : trace_data
`endif
         };
end
`endif

      return output_stage2;

   endfunction

   // -------------------------------------------------------------

   // Initiate DM, Shifter box, MBox or FBox op

   function Action fa_enq (Data_Stage1_to_Stage2 x);
      action
	 rg_stage2  <= x;

	 let funct3 = instr_funct3 (x.instr);

	 // If DMem access, initiate it
`ifdef ISA_A
	 Bool op_stage2_amo = (x.op_stage2 == OP_Stage2_AMO);
	 Bit #(7) amo_funct7 = x.val1 [6:0];
`else
	 Bool op_stage2_amo = False;
	 Bit #(7) amo_funct7 = 0;
`endif
	 if ((x.op_stage2 == OP_Stage2_LD) || (x.op_stage2 == OP_Stage2_ST) || op_stage2_amo) begin
	    WordXL   mstatus     = csr_regfile.read_mstatus;
`ifdef ISA_PRIV_S
	    Bit #(1) sstatus_SUM = (csr_regfile.read_sstatus) [18];
`else
	    Bit #(1) sstatus_SUM = 0;
`endif
	    Bit #(1) mstatus_MXR = mstatus [19];
	    Priv_Mode  mem_priv = x.priv;
	    if (mstatus [17] == 1'b1) begin
	       mem_priv = mstatus [12:11];
	       // $display ("    S2.fa_enq: mem_priv %0d => %0d (mstatus.MPP) due to mstatus.MPRV", x.priv, mem_priv);
	    end

	    CacheOp cache_op = ?;
	    if      (x.op_stage2 == OP_Stage2_LD)  cache_op = CACHE_LD;
	    else if (x.op_stage2 == OP_Stage2_ST)  cache_op = CACHE_ST;
`ifdef ISA_A
	    else if (x.op_stage2 == OP_Stage2_AMO) cache_op = CACHE_AMO;
`endif

            // Prepare the store value
`ifdef RV64
            Bit# (64) wdata_from_gpr = x.val2;
`else
            Bit# (64) wdata_from_gpr = zeroExtend (x.val2);
`endif

`ifdef ISA_F
`ifdef ISA_D
            Bit# (64) wdata_from_fpr = x.fval2;
`else
            Bit# (64) wdata_from_fpr = zeroExtend (x.fval2);
`endif
`ifdef POSIT
            Bit# (64) wdata_from_ppr = zeroExtend (x.pval2);
`endif
`endif
	    dcache.req (cache_op,
			instr_funct3 (x.instr),
`ifdef ISA_A
			amo_funct7,
`endif
			x.addr,
`ifdef ISA_F
`ifdef POSIT
			(x.rs_frm_ppr ? wdata_from_ppr 
                                      : x.rs_frm_fpr ? wdata_from_fpr
                                                     : wdata_from_gpr),
`else
			(x.rs_frm_fpr ? wdata_from_fpr : wdata_from_gpr),
`endif
`else
			wdata_from_gpr,
`endif
			mem_priv,
			sstatus_SUM,
			mstatus_MXR,
			csr_regfile.read_satp);
	 end

`ifdef SHIFT_SERIAL
	 // If Shifter box op, initiate it
	 else if (x.op_stage2 == OP_Stage2_SH)
	    shifter_box.req (unpack (funct3 [2]), x.val1, x.val2);
`endif

`ifdef ISA_M
	 // If MBox op, initiate it
	 else if (x.op_stage2 == OP_Stage2_M) begin
            // Instr fields required for decode for F/D opcodes
	    Bool is_OP_not_OP_32 = (x.instr [3] == 1'b0);
            mbox.req (is_OP_not_OP_32, funct3, x.val1, x.val2);
	 end
`endif

`ifdef ISA_F
	 // If FBox op, initiate it
	 else if (x.op_stage2 == OP_Stage2_FD) begin
	    // Instr fields required for decode for F/D opcodes
            let opcode = instr_opcode (x.instr);
	    let funct7 = instr_funct7 (x.instr);
            let rs2    = instr_rs2    (x.instr);
            Bit #(64) val1 = x.val1_frm_gpr ? extend (x.val1)
                                            : extend (x.fval1);

	    fbox.req (  opcode
		      , funct7
		      , x.rounding_mode   // rm
		      , rs2
		      , val1
		      , extend (x.fval2)
		      , extend (x.fval3) 
`ifdef POSIT
		      , x.pval1
		      , x.pval2 
`endif
		     );
         end
`endif

`ifdef ROCC
	 // If PositAccel op, initiate it
	 else if (x.op_stage2 == OP_Stage2_ROCC) begin
	    // Instr fields required for decode for opcodes
            let opcode = instr_opcode (x.instr);
	    let funct7 = instr_funct7 (x.instr);
            let funct3 = instr_funct3 (x.instr);
            let rs2    = instr_rs2    (x.instr);
            /*Bit #(32) val1 = x.val1_frm_gpr ? extend (x.val1)
                                            : extend (x.fval1);*/ //when dealing with vectors,it maybe used

	    wrap.req (  opcode       //PositAccel is instantiated using wrap
		      , funct7
		      , x.rounding_mode   // rm
		      , funct3          
		      , x.rocc_value_bit           //value bit (RoCC)
                      //,rs2
                      ,x.rd
		      , x.roccval1
		      , x.roccval2
		     );
         end
`endif


`ifdef ACCEL
	 // If PositAccel op, initiate it
	 else if (x.op_stage2 == OP_Stage2_ACCEL) begin
	    // Instr fields required for decode for opcodes
            let opcode = instr_opcode (x.instr);
	    let funct7 = instr_funct7 (x.instr);
            let funct3 = instr_funct3 (x.instr);
            let rs2    = instr_rs2    (x.instr);
            /*Bit #(32) val1 = x.val1_frm_gpr ? extend (x.val1)
                                            : extend (x.fval1);*/ //when dealing with vectors,it maybe used

	    wrap.req (  opcode       //PositAccel is instantiated using wrap
		      , funct7
		      , x.rounding_mode   // rm
		      , funct3          
		      , x.rocc_value_bit           //value bit (RoCC)
                      //,rs2
                      ,x.rd
		      , x.accelval1
		      , x.accelval2
		     );
         end
`endif

      endaction
   endfunction

   // ----------------------------------------------------------------
   // INTERFACE

   // ---- Reset
   interface server_reset = toGPServer (f_reset_reqs, f_reset_rsps);

   // ---- Output
   method Output_Stage2  out;
      return fv_out;
   endmethod

   method Action deq ();
      noAction;
   endmethod

   // ---- Input
   method Action enq (Data_Stage1_to_Stage2 x);
      fa_enq (x);

      if (verbosity > 1)
	 $display ("    CPU_Stage2.enq (Data_Stage1_to_Stage2) ", fshow (x));
   endmethod

   method Action set_full (Bool full);
      rg_full <= full;
   endmethod
endmodule

// ================================================================

endpackage
