// Copyright (c) 2016-2019 Bluespec, Inc. All Rights Reserved

package CPU_Stage1;

// ================================================================
// This is Stage 1 of the "Flute" CPU.
// It contains the EX functionality.
// EX: "Execute"

// ================================================================
// Exports

export
CPU_Stage1_IFC (..),
mkCPU_Stage1;

// ================================================================
// BSV library imports

import FIFOF        :: *;
import GetPut       :: *;
import ClientServer :: *;
import ConfigReg    :: *;

// ----------------
// BSV additional libs

import Cur_Cycle :: *;

// ================================================================
// Project imports

import ISA_Decls        :: *;
import CPU_Globals      :: *;
import Near_Mem_IFC     :: *;
import GPR_RegFile      :: *;
`ifdef ISA_F
import FPR_RegFile      :: *;
`ifdef POSIT
import PPR_RegFile      :: *;
`endif
`endif
`ifdef ACCEL                       //if accelerator is set;assuming both inputs as scalars  and scalar output for now
import PPR_RegFile      :: *;
`endif
import CSR_RegFile      :: *;
import EX_ALU_functions :: *;

`ifdef ISA_C
// 'C' extension (16b compressed instructions)
import CPU_Decode_C     :: *;
`endif

// ================================================================
// Interface

interface CPU_Stage1_IFC;
   // ---- Reset
   interface Server #(Token, Token) server_reset;

   // ---- Output
   (* always_ready *)
   method Output_Stage1 out;

   (* always_ready *)
   method Action deq;

   // ---- Input
   (* always_ready *)
   method Action enq (Data_StageD_to_Stage1  data);

   (* always_ready *)
   method Action set_full (Bool full);
endinterface

// ================================================================
// Implementation module

module mkCPU_Stage1 #(Bit #(4)         verbosity,
		      GPR_RegFile_IFC  gpr_regfile,
		      Bypass           bypass_from_stage2,
		      Bypass           bypass_from_stage3,
`ifdef ISA_F
		      FPR_RegFile_IFC  fpr_regfile,
		      FBypass          fbypass_from_stage2,
		      FBypass          fbypass_from_stage3,
`ifdef POSIT
                      PPR_RegFile_IFC  ppr_regfile,
		      PBypass          pbypass_from_stage2,
		      PBypass          pbypass_from_stage3,
`endif
`endif
`ifdef ACCEL     //asuming that for now dealing with scalars,so just using PPR
                      PPR_RegFile_IFC      ppr_regfile,
		      AccelBypass          accelbypass_from_stage2,
		      AccelBypass          accelbypass_from_stage3,
`endif
		      CSR_RegFile_IFC  csr_regfile,
		      Epoch            cur_epoch,
		      Priv_Mode        cur_priv)
                    (CPU_Stage1_IFC);

   FIFOF #(Token) f_reset_reqs <- mkFIFOF;
   FIFOF #(Token) f_reset_rsps <- mkFIFOF;

   Reg #(Bool)                  rg_full        <- mkReg (False);
   Reg #(Data_StageD_to_Stage1) rg_stage_input <- mkRegU;

   MISA misa   = csr_regfile.read_misa;
   Bit #(2) xl = ((xlen == 32) ? misa_mxl_32 : misa_mxl_64);

   // ----------------------------------------------------------------
   // BEHAVIOR

   rule rl_reset;
      f_reset_reqs.deq;
      rg_full <= False;
      f_reset_rsps.enq (?);
   endrule

   // ----------------
   // ALU

   let decoded_instr  = rg_stage_input.decoded_instr;
   let funct3         = decoded_instr.funct3;
   let funct7         = decoded_instr.funct7;  //func7 of decoded instruction,for the case of accelerator func7 tells which accelerator operation to be performed.

   // Register rs1 read and bypass
   let rs1 = decoded_instr.rs1;
   let rs1_val = gpr_regfile.read_rs1 (rs1);
   match { .busy1a, .rs1a } = fn_gpr_bypass (bypass_from_stage3, rs1, rs1_val);
   match { .busy1b, .rs1b } = fn_gpr_bypass (bypass_from_stage2, rs1, rs1a);
   Bool rs1_busy = (busy1a || busy1b);
   Word rs1_val_bypassed = ((rs1 == 0) ? 0 : rs1b);

   // Register rs2 read and bypass
   let rs2 = decoded_instr.rs2;
   let rs2_val = gpr_regfile.read_rs2 (rs2);
   match { .busy2a, .rs2a } = fn_gpr_bypass (bypass_from_stage3, rs2, rs2_val);
   match { .busy2b, .rs2b } = fn_gpr_bypass (bypass_from_stage2, rs2, rs2a);
   Bool rs2_busy = (busy2a || busy2b);
   Word rs2_val_bypassed = ((rs2 == 0) ? 0 : rs2b);

`ifdef ISA_F
   // FP Register rs1 read and bypass
   let frs1_val = fpr_regfile.read_rs1 (rs1);
   match { .fbusy1a, .frs1a } = fn_fpr_bypass (fbypass_from_stage3, rs1, frs1_val);
   match { .fbusy1b, .frs1b } = fn_fpr_bypass (fbypass_from_stage2, rs1, frs1a);
   Bool frs1_busy = (fbusy1a || fbusy1b);
   WordFL frs1_val_bypassed = frs1b;

   // FP Register rs2 read and bypass
   let frs2_val = fpr_regfile.read_rs2 (rs2);
   match { .fbusy2a, .frs2a } = fn_fpr_bypass (fbypass_from_stage3, rs2, frs2_val);
   match { .fbusy2b, .frs2b } = fn_fpr_bypass (fbypass_from_stage2, rs2, frs2a);
   Bool frs2_busy = (fbusy2a || fbusy2b);
   WordFL frs2_val_bypassed = frs2b;

   // FP Register rs3 read and bypass
   let rs3 = decoded_instr.rs3;
   let frs3_val = fpr_regfile.read_rs3 (rs3);
   match { .fbusy3a, .frs3a } = fn_fpr_bypass (fbypass_from_stage3, rs3, frs3_val);
   match { .fbusy3b, .frs3b } = fn_fpr_bypass (fbypass_from_stage2, rs3, frs3a);
   Bool frs3_busy = (fbusy3a || fbusy3b);
   WordFL frs3_val_bypassed = frs3b;

`ifdef POSIT
   // Posit Register rs1 read and bypass
   let prs1_val = ppr_regfile.read_rs1 (rs1);
   match { .pbusy1a, .prs1a } = fn_ppr_bypass (pbypass_from_stage3, rs1, prs1_val);
   match { .pbusy1b, .prs1b } = fn_ppr_bypass (pbypass_from_stage2, rs1, prs1a);
   Bool prs1_busy = (pbusy1a || pbusy1b);
   WordPL prs1_val_bypassed = prs1b;

   // FP Register rs2 read and bypass
   let prs2_val = ppr_regfile.read_rs2 (rs2);
   match { .pbusy2a, .prs2a } = fn_ppr_bypass (pbypass_from_stage3, rs2, prs2_val);
   match { .pbusy2b, .prs2b } = fn_ppr_bypass (pbypass_from_stage2, rs2, prs2a);
   Bool prs2_busy = (pbusy2a || pbusy2b);
   WordPL prs2_val_bypassed = prs2b;
`endif
`endif

`ifdef ACCEL
   // rs1 read and bypass(similar to POSIT)
   let accelrs1_val = ppr_regfile.read_rs1 (rs1);  
   match { .accelbusy1a, .accelrs1a } = acccel_fn_ppr_bypass (accelbypass_from_stage3, rs1, accelrs1_val);
   match { .accelbusy1b, .accelrs1b } = accel_fn_ppr_bypass (accelbypass_from_stage2, rs1, accelrs1a);
   Bool accelrs1_busy = (accelbusy1a || accelbusy1b);
   WordPL accelrs1_val_bypassed = accelrs1b;

   // rs2 read and bypass(similar to POSIT)
   let accelrs2_val = ppr_regfile.read_rs2 (rs2);
   match { .accelbusy2a, .accelrs2a } = accel_fn_ppr_bypass (pbypass_from_stage3, rs2, accelrs2_val);
   match { .accelbusy2b, .accelrs2b } = accel_fn_ppr_bypass (pbypass_from_stage2, rs2, accelrs2a);
   Bool accelrs2_busy = (accelbusy2a || accelbusy2b);
   WordPL accelrs2_val_bypassed = accelrs2b;
`endif


   // ALU function
   let alu_inputs = ALU_Inputs {cur_priv       : cur_priv,
				pc             : rg_stage_input.pc,
				is_i32_not_i16 : rg_stage_input.is_i32_not_i16,
				instr          : rg_stage_input.instr,//32 bit instruction 
`ifdef ISA_C
				instr_C        : rg_stage_input.instr_C,
`endif
				decoded_instr  : rg_stage_input.decoded_instr,//decoded instruction
				rs1_val        : rs1_val_bypassed,
				rs2_val        : rs2_val_bypassed,
`ifdef ISA_F
				frs1_val       : frs1_val_bypassed,
				frs2_val       : frs2_val_bypassed,
				frs3_val       : frs3_val_bypassed,
				frm            : csr_regfile.read_frm,
`ifdef INCLUDE_TANDEM_VERIF
                                fflags         : csr_regfile.read_fflags,
`endif

`ifdef POSIT
				prs1_val       : prs1_val_bypassed,
				prs2_val       : prs2_val_bypassed,
`endif
`endif

`ifdef ACCEL 
				accelrs1_val   : accelrs1_val_bypassed,
				accelrs2_val   : accelrs2_val_bypassed,
				rocc_value_bit : rg_stage_input.rocc_value_bit,  //value bit of RoCC
`endif
				mstatus        : csr_regfile.read_mstatus,
				misa           : csr_regfile.read_misa };

   let alu_outputs = fv_ALU (alu_inputs);

   let data_to_stage2 = Data_Stage1_to_Stage2 {pc            : rg_stage_input.pc,
					       instr         : rg_stage_input.instr,
					       op_stage2     : alu_outputs.op_stage2,
					       rd            : alu_outputs.rd,
					       addr          : alu_outputs.addr,
					       val1          : alu_outputs.val1,
					       val2          : alu_outputs.val2,
`ifdef ISA_F
					       fval1         : alu_outputs.fval1,
					       fval2         : alu_outputs.fval2,
					       fval3         : alu_outputs.fval3,
					       rd_in_fpr     : alu_outputs.rd_in_fpr,
					       rs_frm_fpr    : alu_outputs.rs_frm_fpr,
					       val1_frm_gpr  : alu_outputs.val1_frm_gpr,
`ifdef POSIT
                           no_rd_upd     : alu_outputs.no_rd_upd,
					       rs_frm_ppr    : alu_outputs.rs_frm_ppr,
					       rd_in_ppr     : alu_outputs.rd_in_ppr,
					       pval1         : alu_outputs.pval1,
					       pval2         : alu_outputs.pval2,
`endif
					       rounding_mode : alu_outputs.rm,
`endif

`ifdef ACCEL            //ToDo:include GPR when dealing with vectors
                          
					       accelval1     : alu_outputs.accelval1,//input1
					       accelval2     : alu_outputs.accelval2,//input2
						   rs_frm_ppr    : alu_outputs.rs_frm_ppr,
					       rd_in_ppr     : alu_outputs.rd_in_ppr,
						   funct3        : alu_outputs.funct3, //In RoCC,funct3 is referred as rg_sel=[xd xs1 xs2]
                           no_rd_upd     : alu_outputs.no_rd_upd,
						   funct7	     : alu_outputs.funct7, //in accelerator funct7 acts as the opcode to determine what accelerator operation to be carried out
						   rocc_value_bit : alu_outputs.rocc_value_bit,  //value bit for RoCC
						   rounding_mode : alu_outputs.rm,
`endif
`ifdef INCLUDE_TANDEM_VERIF
					       trace_data    : alu_outputs.trace_data,
`endif
					       priv          : cur_priv };

   // ----------------
   // Combinational output function

   function Output_Stage1 fv_out;
      Output_Stage1 output_stage1 = ?;

      // This stage is empty
      if (! rg_full) begin
	 output_stage1.ostatus = OSTATUS_EMPTY;
      end

      // Wrong branch-prediction epoch: discard instruction (convert into a NOOP)
      else if (rg_stage_input.epoch != cur_epoch) begin
	 output_stage1.ostatus = OSTATUS_PIPE;
	 output_stage1.control = CONTROL_DISCARD;

	 // For debugging only
	 let data_to_stage2 = Data_Stage1_to_Stage2 {pc:        rg_stage_input.pc,
						     instr:     rg_stage_input.instr,
						     op_stage2: OP_Stage2_ALU,
						     rd:        0,
						     addr:      ?,
						     val1:      ?,
						     val2:      ?,
`ifdef ISA_F
						     fval1           : ?,
						     fval2           : ?,
						     fval3           : ?,
						     rd_in_fpr       : ?,
					         rs_frm_fpr      : ?,
					         val1_frm_gpr    : ?,
`ifdef POSIT
						     pval1           : ?,
						     pval2           : ?,
					         rs_frm_ppr      : ?,
						     rd_in_ppr       : ?,
                             no_rd_upd       : ?,
`endif
						     rounding_mode   : ?,
`endif

`ifdef ACCEL
						     accelval1           : ?,
						     accelval2           : ?,
					         rs_frm_ppr      : ?,
						     rd_in_ppr       : ?,
							 no_rd_upd       : ?,
                             funct3          : ?,
                             funct7		     : ?,
							 rocc_value_bit  : ?,
							 rounding_mode   : ?,
							
`endif


`ifdef INCLUDE_TANDEM_VERIF
						     trace_data: alu_outputs.trace_data,
`endif
						     priv:      cur_priv
						     };

	 output_stage1.data_to_stage2 = data_to_stage2;
      end

      // Stall if bypass pending for GPR rs1 or rs2
      else if (rs1_busy || rs2_busy) begin
	 output_stage1.ostatus = OSTATUS_BUSY;
      end

`ifdef ISA_F
      // Stall if bypass pending for FPR rs1, rs2 or rs3
      else if (frs1_busy || frs2_busy || frs3_busy) begin
	 output_stage1.ostatus = OSTATUS_BUSY;
      end
`ifdef POSIT
      // Stall if bypass pending for PPR rs1, rs2 or rs3
      else if (prs1_busy || prs2_busy) begin
	 output_stage1.ostatus = OSTATUS_BUSY;
      end
`endif
`endif
`ifdef ACCEL
      // Stall if bypass pending for PPR rs1, rs2 or rs3
      else if (accelrs1_busy || accelrs2_busy) begin
	 output_stage1.ostatus = OSTATUS_BUSY;
      end
`endif

      // Trap on fetch-exception
      else if (rg_stage_input.exc) begin
	 output_stage1.ostatus   = OSTATUS_NONPIPE;
	 output_stage1.control   = CONTROL_TRAP;
	 output_stage1.trap_info = Trap_Info {epc:      rg_stage_input.pc,
					      exc_code: rg_stage_input.exc_code,
					      tval:     rg_stage_input.tval};
	 output_stage1.data_to_stage2 = data_to_stage2;
      end

      // ALU outputs: pipe (straight/branch)
      // and non-pipe (CSRR_W, CSRR_S_or_C, FENCE.I, FENCE, SFENCE_VMA, xRET, WFI, TRAP)
      else begin
	 let ostatus = (  (   (alu_outputs.control == CONTROL_STRAIGHT)
			   || (alu_outputs.control == CONTROL_BRANCH))
			? OSTATUS_PIPE
			: OSTATUS_NONPIPE);

	 // Compute MTVAL in case of traps
	 let tval = 0;
	 if (alu_outputs.exc_code == exc_code_ILLEGAL_INSTRUCTION) begin
	    // The instruction
`ifdef ISA_C
	    tval = (rg_stage_input.is_i32_not_i16
		    ? zeroExtend (rg_stage_input.instr)
		    : zeroExtend (rg_stage_input.instr_C));
`else
	    tval = zeroExtend (rg_stage_input.instr);
`endif
	 end
	 else if (alu_outputs.exc_code == exc_code_INSTR_ADDR_MISALIGNED)
	    tval = alu_outputs.addr;                           // The branch target pc
	 else if (alu_outputs.exc_code == exc_code_BREAKPOINT)
	    tval = rg_stage_input.pc;                          // The faulting virtual address

	 let trap_info = Trap_Info {epc:      rg_stage_input.pc,
				    exc_code: alu_outputs.exc_code,
				    tval:     tval};

	 let fall_through_pc = rg_stage_input.pc + (rg_stage_input.is_i32_not_i16 ? 4 : 2);
	 let next_pc = ((alu_outputs.control == CONTROL_BRANCH)
			? alu_outputs.addr
			: fall_through_pc);
	 let redirect = (next_pc != rg_stage_input.pred_pc);

	 output_stage1.ostatus        = ostatus;
	 output_stage1.control        = alu_outputs.control;
	 output_stage1.trap_info      = trap_info;
	 output_stage1.redirect       = redirect;
	 output_stage1.next_pc        = next_pc;
	 output_stage1.cf_info        = alu_outputs.cf_info;
	 output_stage1.data_to_stage2 = data_to_stage2;
      end

      return output_stage1;
   endfunction: fv_out

   // ================================================================
   // INTERFACE

   // ---- Reset
   interface server_reset = toGPServer (f_reset_reqs, f_reset_rsps);

   // ---- Output
   method Output_Stage1 out;
      return fv_out;
   endmethod

   method Action deq ();
   endmethod

   // ---- Input
   method Action enq (Data_StageD_to_Stage1  data);
      rg_stage_input <= data;
      if (verbosity > 1)
	 $display ("    CPU_Stage1.enq: 0x%08h", data.pc);
   endmethod

   method Action set_full (Bool full);
      rg_full <= full;
   endmethod
endmodule

// ================================================================

endpackage
